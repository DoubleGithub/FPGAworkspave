LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL; 
ENTITY CNT4B_S IS
PORT (CLK : IN STD_LOGIC;
      CQ : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
      CQ_DELAY : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END CNT4B_S;
ARCHITECTURE behav OF CNT4B_S IS 
SIGNAL CQI : STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
PROCESS(CLK)
BEGIN
 IF CLK'EVENT AND CLK='1' THEN
    CQI <= CQI + 1;	
    CQ_DELAY <= CQI  ; 
 END IF; 
 CQ <= CQI;
END PROCESS;
END behav;