LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL; 
ENTITY SCAN_LED IS
PORT ( CLK : IN STD_LOGIC; 
LK   : IN STD_LOGIC;
DIN	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
DP  : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
SG	: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);  --�ο����ź����
BT	: OUT STD_LOGIC_VECTOR(7 DOWNTO 0) );--λ�����ź����
END;
ARCHITECTURE one OF SCAN_LED IS
SIGNAL CNT8  : STD_LOGIC_VECTOR(2 DOWNTO 0); 
SIGNAL DOUT  : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	A  : STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
P1:PROCESS( LK,DIN)
BEGIN
IF LK'EVENT	AND LK	= '1'THEN DOUT <= DIN; 
END IF;
END PROCESS P1;
P2:PROCESS( CNT8 )
BEGIN
CASE  CNT8  IS
WHEN "000" =>  BT <= "11111110" ; A <= DOUT(3 DOWNTO 0) ; SG(7) <= DP(0);
WHEN "001" =>  BT <= "11111101" ; A <= DOUT(7 DOWNTO 4) ; SG(7) <= DP(1);
WHEN "010" =>  BT <= "11111011" ; A <= DOUT(11 DOWNTO 8) ; SG(7) <= DP(2);
WHEN "011" =>  BT <= "11110111" ; A <= DOUT(15 DOWNTO 12) ; SG(7) <= DP(3);
WHEN "100" =>  BT <= "11101111" ; A <= DOUT(19 DOWNTO 16) ; SG(7) <= DP(4);
WHEN "101" =>  BT <= "11011111" ; A <= DOUT(23 DOWNTO 20) ; SG(7) <= DP(5);
WHEN "110" =>  BT <= "10111111" ; A <= DOUT(27 DOWNTO 24) ; SG(7) <= DP(6);
WHEN "111" =>  BT <= "01111111" ; A <= DOUT(31 DOWNTO 28) ; SG(7) <= DP(7);
WHEN OTHERS =>  NULL ;
END CASE ;
END PROCESS P2;
P3:PROCESS(CLK)
BEGIN
IF CLK'EVENT AND CLK = '1' THEN 
CNT8 <= CNT8 + 1; 
END IF;
END PROCESS P3; 
P4:PROCESS( A ) --�����·
BEGIN 
CASE  A  IS
WHEN "0000"	=> SG(6 DOWNTO 0) <= "0111111";  WHEN "0001" => SG(6 DOWNTO 0) <= "0000110";
WHEN "0010"	=> SG(6 DOWNTO 0) <= "1011011";  WHEN "0011" => SG(6 DOWNTO 0) <= "1001111";
WHEN "0100"	=> SG(6 DOWNTO 0) <= "1100110";  WHEN "0101" => SG(6 DOWNTO 0) <= "1101101";
WHEN "0110"	=> SG(6 DOWNTO 0) <= "1111101";  WHEN "0111" => SG(6 DOWNTO 0) <= "0000111";
WHEN "1000"	=> SG(6 DOWNTO 0) <= "1111111";  WHEN "1001" => SG(6 DOWNTO 0) <= "1101111";
WHEN "1010" => SG(6 DOWNTO 0) <= "1110111";  WHEN "1011" => SG(6 DOWNTO 0) <= "1111100"; 
WHEN "1100" => SG(6 DOWNTO 0) <= "0111001";  WHEN "1101" => SG(6 DOWNTO 0) <= "1011110"; 
WHEN "1110" => SG(6 DOWNTO 0) <= "1111001";  WHEN "1111" => SG(6 DOWNTO 0) <= "1110001"; 
WHEN OTHERS =>  NULL ;
END CASE ;
END PROCESS P4; 
END;
