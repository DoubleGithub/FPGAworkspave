LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL; 
ENTITY data_bus IS
PORT (CLK : IN STD_LOGIC;
            
      ----M[3..0]=0001
      SW : OUT STD_LOGIC_VECTOR(16 DOWNTO 1);
      
      ----M[3..0]=0011
      PB : OUT STD_LOGIC_VECTOR(16 DOWNTO 1);
      
      ----M[3..0]=0111
      LED : IN STD_LOGIC_VECTOR(16 DOWNTO 1);
      
      ----M[3..0]=0010
      SEG : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      COM : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      
      ----M[3..0]=0101
      ROW : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
      COL : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      
      ----M[3..0]=0110
      DOT : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
      ADDRESS : IN STD_LOGIC_VECTOR(4 DOWNTO 1);
      
      ----------------------------------------------
      Mout : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
      D : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
      A : OUT STD_LOGIC_VECTOR(4 DOWNTO 1));
END;
ARCHITECTURE behav OF data_bus IS
 SIGNAL Mtemp : STD_LOGIC_VECTOR(3 DOWNTO 0);
 SIGNAL CQI : STD_LOGIC_VECTOR(2 DOWNTO 0);
 SIGNAL SWtemp,PBtemp : STD_LOGIC_VECTOR(16 DOWNTO 1);
 SIGNAL ROWtemp : STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
 Mout <= Mtemp;
 PROCESS(CLK)
BEGIN
 IF CLK'EVENT AND CLK='1' THEN
  IF CQI < 5 THEN
    CQI <= CQI + 1;
  ELSE	
    CQI <= "000"; 
 END IF; 
 END IF;
END PROCESS;
PROCESS(CQI)
BEGIN
 CASE CQI IS
 WHEN "000" => Mtemp<="0001";
 WHEN "001" => Mtemp<="0011";
 WHEN "010" => Mtemp<="0111";
 WHEN "011" => Mtemp<="0010";
 WHEN "100" => Mtemp<="0101";
 WHEN "101" => Mtemp<="0110";
 WHEN OTHERS => NULL;
 END CASE;
END PROCESS;
 
 PROCESS(CLK,Mtemp,LED,SEG,COM,COL,DOT,ADDRESS,D)
 BEGIN
 
  CASE Mtemp IS
  WHEN "0001" => SWtemp(16 DOWNTO 1)<=D(15 DOWNTO 0);D<=(OTHERS=>'Z');
  WHEN "0011" => PBtemp(16 DOWNTO 1)<=D(15 DOWNTO 0);D<=(OTHERS=>'Z');
  WHEN "0111" => D(15 DOWNTO 0)<=LED(16 DOWNTO 1);
  WHEN "0010" => D(15 DOWNTO 8) <= COM; D(7 DOWNTO 0) <=SEG;
  WHEN "0101" => D(7 DOWNTO 4)<=COL;D(15 DOWNTO 8)<=(OTHERS=>'Z');D(3 DOWNTO 0)<=(OTHERS=>'Z');ROWtemp<=D(3 DOWNTO 0);             
  WHEN "0110" => D <= DOT;A<=ADDRESS;
  WHEN OTHERS => D<=(OTHERS=>'Z');
  END CASE;
  IF CLK'EVENT AND CLK='0' THEN
   SW <=SWtemp;
   PB <=PBtemp;
   ROW <=ROWtemp;
  END IF;
 END PROCESS;
END;