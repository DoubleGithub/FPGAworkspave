LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL; 

ENTITY sikaoti IS
PORT (CLK : IN STD_LOGIC;
      RST,EN,LD : IN STD_LOGIC;
      DIN : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
      CQ : OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
END sikaoti;
ARCHITECTURE behav OF sikaoti IS
BEGIN
PROCESS(CLK, RST, EN)
 VARIABLE CQI : STD_LOGIC_VECTOR(4 DOWNTO 0):= B"11000";
BEGIN
 IF RST = '1' THEN	
    --CQI := (OTHERS =>'0') ;
    CQI := B"11000" ;
 ELSIF CLK'EVENT AND CLK='1' THEN	
    IF LD = '1' THEN
       CQI := DIN;
    ELSIF EN = '1' THEN
       CQI := CQI - 1;
    END IF;
 END IF; 

 IF CQI = 0 THEN 
    CQI := B"11000" ;  
 END IF;
 CQ <= CQI;
END PROCESS;
END behav;