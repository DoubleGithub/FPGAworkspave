LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL; 
ENTITY CNT4B IS
PORT (CLK : IN STD_LOGIC;
      RST,EN,LD : IN STD_LOGIC;
      DIN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      CQ : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
      COUT : OUT STD_LOGIC);
END CNT4B;
ARCHITECTURE behav OF CNT4B IS
BEGIN
PROCESS(CLK, RST, EN)
 VARIABLE CQI : STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
 IF RST = '1' THEN	
    CQI := (OTHERS =>'0') ;
 ELSIF CLK'EVENT AND CLK='1' THEN	
    IF LD = '1' THEN
       CQI := DIN;
    ELSIF EN = '1' THEN
       CQI := CQI + 1;
    END IF;
 END IF; 

 IF CQI = 15 THEN 
    COUT <= '1';
 ELSE 
    COUT <= '0'; 
 END IF;
 CQ <= CQI;
END PROCESS;
END behav;